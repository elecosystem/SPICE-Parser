*Simple linear example

example exercise
V1 1 0 2V
R1 1 2 2ohm
Vm 2 3 0V;
V2 1 0 Vm 2
R2 3 0 2V
.END
